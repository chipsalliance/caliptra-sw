// SPDX-License-Identifier: Apache-2.0
// Stub module for AXI4 Protocol Checker - not needed for verilator simulation

// Empty module - AXI4PC is not synthesized in verilator
module Axi4PC;
endmodule
